----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04.04.2024 13:55:04
-- Design Name: 
-- Module Name: comparator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

-- Programa para comparar
entity comparator is

    Port ( A : in unsigned(4 downto 0);
           B : in unsigned(4 downto 0);
           equal : out std_logic);
end comparator;

architecture Behavioral of comparator is

begin
    Process(A,B)
        begin
            if A = B then
                    equal <= '1';
                else
                equal <= '0'; 
            end if;               
    end process;
end Behavioral;
